<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>42.4932,-31.4674,205.694,-112.134</PageViewport>
<gate>
<ID>1</ID>
<type>GA_LED</type>
<position>94,-101.5</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>52,-41</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>3</ID>
<type>GA_LED</type>
<position>74.5,-40.5</position>
<input>
<ID>N_in0</ID>3 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>4</ID>
<type>AA_LABEL</type>
<position>45.5,-40.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>5</ID>
<type>AA_LABEL</type>
<position>81.5,-40</position>
<gparam>LABEL_TEXT Output Y=A'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>6</ID>
<type>AA_LABEL</type>
<position>66,-33.5</position>
<gparam>LABEL_TEXT NOR as NOT Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>7</ID>
<type>AA_LABEL</type>
<position>101,-101</position>
<gparam>LABEL_TEXT Output Y=(A.B)'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>GA_LED</type>
<position>81.5,-56.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>9</ID>
<type>AA_LABEL</type>
<position>88.5,-56</position>
<gparam>LABEL_TEXT Output Y=A+B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_TOGGLE</type>
<position>50,-55.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>43.5,-55</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_TOGGLE</type>
<position>50,-58.5</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>13</ID>
<type>BE_NOR2</type>
<position>63.5,-40.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>44,-58.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>66,-50</position>
<gparam>LABEL_TEXT NOR as OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>85.5,-77</position>
<input>
<ID>N_in0</ID>14 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>BE_NOR2</type>
<position>59.5,-57</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>92.5,-76.5</position>
<gparam>LABEL_TEXT Output Y=A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>19</ID>
<type>BE_NOR2</type>
<position>73,-57</position>
<input>
<ID>IN_0</ID>7 </input>
<input>
<ID>IN_1</ID>7 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>53,-73.5</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_LABEL</type>
<position>46.5,-73</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_TOGGLE</type>
<position>53,-82</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>47.5,-82</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>70,-66.5</position>
<gparam>LABEL_TEXT NOR as AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_TOGGLE</type>
<position>54,-97</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>47.5,-96.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>BE_NOR2</type>
<position>62.5,-73.5</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>AA_TOGGLE</type>
<position>54,-105.5</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>29</ID>
<type>BE_NOR2</type>
<position>62.5,-82</position>
<input>
<ID>IN_0</ID>15 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>48.5,-105.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>BE_NOR2</type>
<position>75.5,-78</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>71,-90</position>
<gparam>LABEL_TEXT NOR as NAND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>BE_NOR2</type>
<position>63.5,-97</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>34</ID>
<type>BE_NOR2</type>
<position>63.5,-105.5</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>35</ID>
<type>BE_NOR2</type>
<position>76.5,-101.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>17 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>36</ID>
<type>GA_LED</type>
<position>173,-39</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>BE_NOR2</type>
<position>85.5,-101.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>AA_LABEL</type>
<position>182,-38.5</position>
<gparam>LABEL_TEXT Output Y=A'B+AB'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>39</ID>
<type>AA_TOGGLE</type>
<position>130.5,-35.5</position>
<output>
<ID>OUT_0</ID>27 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_LABEL</type>
<position>124,-35</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_TOGGLE</type>
<position>130.5,-44</position>
<output>
<ID>OUT_0</ID>26 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>42</ID>
<type>AA_LABEL</type>
<position>125,-44</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>147.5,-28.5</position>
<gparam>LABEL_TEXT NAND as XOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>50</ID>
<type>BE_NOR2</type>
<position>142,-39.5</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>BE_NOR2</type>
<position>153,-36</position>
<input>
<ID>IN_0</ID>27 </input>
<input>
<ID>IN_1</ID>28 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>54</ID>
<type>BE_NOR2</type>
<position>153,-44.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>26 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>BE_NOR2</type>
<position>160,-40</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>58</ID>
<type>BE_NOR2</type>
<position>167,-40</position>
<input>
<ID>IN_0</ID>32 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>187.5,-70.5</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>196.5,-70</position>
<gparam>LABEL_TEXT Output Y=AB+A'B'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_TOGGLE</type>
<position>128,-66</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>121.5,-65.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_TOGGLE</type>
<position>128,-74.5</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>122.5,-74.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>145,-59</position>
<gparam>LABEL_TEXT NAND as XNOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>BE_NOR2</type>
<position>139.5,-70</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>67</ID>
<type>BE_NOR2</type>
<position>150.5,-66.5</position>
<input>
<ID>IN_0</ID>35 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>68</ID>
<type>BE_NOR2</type>
<position>150.5,-75</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>34 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>69</ID>
<type>BE_NOR2</type>
<position>157.5,-70.5</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>39 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>70</ID>
<type>BE_NOR2</type>
<position>164.5,-70.5</position>
<input>
<ID>IN_0</ID>39 </input>
<input>
<ID>IN_1</ID>39 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>BE_NOR2</type>
<position>174,-70.5</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>AA_LABEL</type>
<position>102.5,-18.5</position>
<gparam>LABEL_TEXT NOR as UNIVERSAL GATES</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-100.5,70,-97</points>
<intersection>-100.5 1</intersection>
<intersection>-97 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-100.5,73.5,-100.5</points>
<connection>
<GID>35</GID>
<name>IN_0</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66.5,-97,70,-97</points>
<connection>
<GID>33</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-105.5,70,-102.5</points>
<intersection>-105.5 2</intersection>
<intersection>-102.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>70,-102.5,73.5,-102.5</points>
<connection>
<GID>35</GID>
<name>IN_1</name></connection>
<intersection>70 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>66.5,-105.5,70,-105.5</points>
<connection>
<GID>34</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>66.5,-40.5,73.5,-40.5</points>
<connection>
<GID>3</GID>
<name>N_in0</name></connection>
<connection>
<GID>13</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-41.5,60.5,-39.5</points>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-41,60.5,-41</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-106.5,60.5,-104.5</points>
<connection>
<GID>34</GID>
<name>IN_1</name></connection>
<connection>
<GID>34</GID>
<name>IN_0</name></connection>
<intersection>-105.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-105.5,60.5,-105.5</points>
<connection>
<GID>28</GID>
<name>OUT_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>70,-58,70,-56</points>
<connection>
<GID>19</GID>
<name>IN_0</name></connection>
<connection>
<GID>19</GID>
<name>IN_1</name></connection>
<intersection>-57 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>62.5,-57,70,-57</points>
<connection>
<GID>17</GID>
<name>OUT</name></connection>
<intersection>70 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>78,-57,78,-56.5</points>
<intersection>-57 2</intersection>
<intersection>-56.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>78,-56.5,80.5,-56.5</points>
<connection>
<GID>8</GID>
<name>N_in0</name></connection>
<intersection>78 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>76,-57,78,-57</points>
<connection>
<GID>19</GID>
<name>OUT</name></connection>
<intersection>78 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-58.5,54,-58</points>
<intersection>-58.5 2</intersection>
<intersection>-58 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-58,56.5,-58</points>
<connection>
<GID>17</GID>
<name>IN_1</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-58.5,54,-58.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>54,-56,54,-55.5</points>
<intersection>-56 1</intersection>
<intersection>-55.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>54,-56,56.5,-56</points>
<connection>
<GID>17</GID>
<name>IN_0</name></connection>
<intersection>54 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-55.5,54,-55.5</points>
<connection>
<GID>10</GID>
<name>OUT_0</name></connection>
<intersection>54 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60.5,-98,60.5,-96</points>
<connection>
<GID>33</GID>
<name>IN_1</name></connection>
<connection>
<GID>33</GID>
<name>IN_0</name></connection>
<intersection>-97 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-97,60.5,-97</points>
<connection>
<GID>25</GID>
<name>OUT_0</name></connection>
<intersection>60.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-77,69,-73.5</points>
<intersection>-77 1</intersection>
<intersection>-73.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-77,72.5,-77</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-73.5,69,-73.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-82,69,-79</points>
<intersection>-82 2</intersection>
<intersection>-79 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-79,72.5,-79</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>65.5,-82,69,-82</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81.5,-78,81.5,-77</points>
<intersection>-78 2</intersection>
<intersection>-77 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>81.5,-77,84.5,-77</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<intersection>81.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>78.5,-78,81.5,-78</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<intersection>81.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-83,59.5,-81</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-82,59.5,-82</points>
<connection>
<GID>22</GID>
<name>OUT_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>59.5,-74.5,59.5,-72.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-73.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-73.5,59.5,-73.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>59.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>81,-102.5,81,-100.5</points>
<intersection>-102.5 2</intersection>
<intersection>-101.5 1</intersection>
<intersection>-100.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>79.5,-101.5,81,-101.5</points>
<connection>
<GID>35</GID>
<name>OUT</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>81,-102.5,82.5,-102.5</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>81 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>81,-100.5,82.5,-100.5</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>81 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>88.5,-101.5,93,-101.5</points>
<connection>
<GID>1</GID>
<name>N_in0</name></connection>
<connection>
<GID>37</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>171,-40,171,-39</points>
<intersection>-40 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>171,-39,172,-39</points>
<connection>
<GID>36</GID>
<name>N_in0</name></connection>
<intersection>171 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>170,-40,171,-40</points>
<connection>
<GID>58</GID>
<name>OUT</name></connection>
<intersection>171 0</intersection></hsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>135.5,-45.5,135.5,-44</points>
<intersection>-45.5 1</intersection>
<intersection>-44 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>135.5,-45.5,150,-45.5</points>
<connection>
<GID>54</GID>
<name>IN_1</name></connection>
<intersection>135.5 0</intersection>
<intersection>139 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>132.5,-44,135.5,-44</points>
<connection>
<GID>41</GID>
<name>OUT_0</name></connection>
<intersection>135.5 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>139,-45.5,139,-40.5</points>
<connection>
<GID>50</GID>
<name>IN_1</name></connection>
<intersection>-45.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>132.5,-35.5,150,-35.5</points>
<connection>
<GID>39</GID>
<name>OUT_0</name></connection>
<intersection>139 4</intersection>
<intersection>150 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>150,-35.5,150,-35</points>
<connection>
<GID>52</GID>
<name>IN_0</name></connection>
<intersection>-35.5 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>139,-38.5,139,-35.5</points>
<connection>
<GID>50</GID>
<name>IN_0</name></connection>
<intersection>-35.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>147.5,-43.5,147.5,-37</points>
<intersection>-43.5 3</intersection>
<intersection>-39.5 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>145,-39.5,147.5,-39.5</points>
<connection>
<GID>50</GID>
<name>OUT</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>147.5,-37,150,-37</points>
<connection>
<GID>52</GID>
<name>IN_1</name></connection>
<intersection>147.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>147.5,-43.5,150,-43.5</points>
<connection>
<GID>54</GID>
<name>IN_0</name></connection>
<intersection>147.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-39,156.5,-36</points>
<intersection>-39 1</intersection>
<intersection>-36 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-39,157,-39</points>
<connection>
<GID>56</GID>
<name>IN_0</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156,-36,156.5,-36</points>
<connection>
<GID>52</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>156.5,-44.5,156.5,-41</points>
<intersection>-44.5 2</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>156.5,-41,157,-41</points>
<connection>
<GID>56</GID>
<name>IN_1</name></connection>
<intersection>156.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>156,-44.5,156.5,-44.5</points>
<connection>
<GID>54</GID>
<name>OUT</name></connection>
<intersection>156.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-41,163.5,-39</points>
<intersection>-41 3</intersection>
<intersection>-40 2</intersection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>163.5,-39,164,-39</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>163,-40,163.5,-40</points>
<connection>
<GID>56</GID>
<name>OUT</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>163.5,-41,164,-41</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>133,-76,133,-74.5</points>
<intersection>-76 1</intersection>
<intersection>-74.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>133,-76,147.5,-76</points>
<connection>
<GID>68</GID>
<name>IN_1</name></connection>
<intersection>133 0</intersection>
<intersection>136.5 4</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>130,-74.5,133,-74.5</points>
<connection>
<GID>63</GID>
<name>OUT_0</name></connection>
<intersection>133 0</intersection></hsegment>
<vsegment>
<ID>4</ID>
<points>136.5,-76,136.5,-71</points>
<connection>
<GID>66</GID>
<name>IN_1</name></connection>
<intersection>-76 1</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>130,-66,147.5,-66</points>
<connection>
<GID>61</GID>
<name>OUT_0</name></connection>
<intersection>136.5 4</intersection>
<intersection>147.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>147.5,-66,147.5,-65.5</points>
<connection>
<GID>67</GID>
<name>IN_0</name></connection>
<intersection>-66 1</intersection></vsegment>
<vsegment>
<ID>4</ID>
<points>136.5,-69,136.5,-66</points>
<connection>
<GID>66</GID>
<name>IN_0</name></connection>
<intersection>-66 1</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>145,-74,145,-67.5</points>
<intersection>-74 3</intersection>
<intersection>-70 1</intersection>
<intersection>-67.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>142.5,-70,145,-70</points>
<connection>
<GID>66</GID>
<name>OUT</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>145,-67.5,147.5,-67.5</points>
<connection>
<GID>67</GID>
<name>IN_1</name></connection>
<intersection>145 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>145,-74,147.5,-74</points>
<connection>
<GID>68</GID>
<name>IN_0</name></connection>
<intersection>145 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-69.5,154,-66.5</points>
<intersection>-69.5 1</intersection>
<intersection>-66.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-69.5,154.5,-69.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>153.5,-66.5,154,-66.5</points>
<connection>
<GID>67</GID>
<name>OUT</name></connection>
<intersection>154 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>154,-75,154,-71.5</points>
<intersection>-75 2</intersection>
<intersection>-71.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>154,-71.5,154.5,-71.5</points>
<connection>
<GID>69</GID>
<name>IN_1</name></connection>
<intersection>154 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>153.5,-75,154,-75</points>
<connection>
<GID>68</GID>
<name>OUT</name></connection>
<intersection>154 0</intersection></hsegment></shape></wire>
<wire>
<ID>39</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>161,-71.5,161,-69.5</points>
<intersection>-71.5 3</intersection>
<intersection>-70.5 2</intersection>
<intersection>-69.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>161,-69.5,161.5,-69.5</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>160.5,-70.5,161,-70.5</points>
<connection>
<GID>69</GID>
<name>OUT</name></connection>
<intersection>161 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>161,-71.5,161.5,-71.5</points>
<connection>
<GID>70</GID>
<name>IN_1</name></connection>
<intersection>161 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>167.5,-70.5,171,-70.5</points>
<connection>
<GID>70</GID>
<name>OUT</name></connection>
<intersection>171 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>171,-71.5,171,-69.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>-70.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>177,-70.5,186.5,-70.5</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>72</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 9></circuit>
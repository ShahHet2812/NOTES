<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>111.574,-13.453,274.775,-94.1202</PageViewport>
<gate>
<ID>51</ID>
<type>AA_LABEL</type>
<position>99,-31.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>52</ID>
<type>AA_LABEL</type>
<position>99,-38.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_TOGGLE</type>
<position>102.5,-32</position>
<output>
<ID>OUT_0</ID>14 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>102,-39</position>
<output>
<ID>OUT_0</ID>15 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>55</ID>
<type>AI_XOR2</type>
<position>112.5,-35.5</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>16 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>56</ID>
<type>GA_LED</type>
<position>118,-35.5</position>
<input>
<ID>N_in0</ID>16 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>57</ID>
<type>AA_INVERTER</type>
<position>111,-45</position>
<input>
<ID>IN_0</ID>14 </input>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>58</ID>
<type>AA_AND2</type>
<position>118,-50.5</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>15 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>59</ID>
<type>GA_LED</type>
<position>125.5,-50.5</position>
<input>
<ID>N_in0</ID>18 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>60</ID>
<type>AA_LABEL</type>
<position>128.5,-35</position>
<gparam>LABEL_TEXT DIFFERENCE(A'B+AB')</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>61</ID>
<type>AA_LABEL</type>
<position>132.5,-50.5</position>
<gparam>LABEL_TEXT BORROW(A'B)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>62</ID>
<type>AA_LABEL</type>
<position>134.5,-18</position>
<gparam>LABEL_TEXT HALF SUBTRACTOR</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>63</ID>
<type>AA_LABEL</type>
<position>174.5,-26</position>
<gparam>LABEL_TEXT AOI</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>64</ID>
<type>AA_LABEL</type>
<position>116,-26</position>
<gparam>LABEL_TEXT SIMPLIFIED DIAGRAM</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>163.5,-30.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_LABEL</type>
<position>174.5,-30.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>67</ID>
<type>AA_TOGGLE</type>
<position>163.5,-35</position>
<output>
<ID>OUT_0</ID>19 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>175,-35</position>
<output>
<ID>OUT_0</ID>20 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_INVERTER</type>
<position>170,-44.5</position>
<input>
<ID>IN_0</ID>19 </input>
<output>
<ID>OUT_0</ID>21 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>70</ID>
<type>AA_INVERTER</type>
<position>183.5,-44</position>
<input>
<ID>IN_0</ID>20 </input>
<output>
<ID>OUT_0</ID>22 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>71</ID>
<type>AA_AND2</type>
<position>193,-54</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>23 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>AA_AND2</type>
<position>193.5,-63</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>24 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>AE_OR2</type>
<position>203,-58.5</position>
<input>
<ID>IN_0</ID>23 </input>
<input>
<ID>IN_1</ID>24 </input>
<output>
<ID>OUT</ID>25 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>GA_LED</type>
<position>207,-58.5</position>
<input>
<ID>N_in0</ID>25 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>75</ID>
<type>AA_LABEL</type>
<position>218,-58.5</position>
<gparam>LABEL_TEXT DIFFERENCE(A'B+AB')</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>76</ID>
<type>AA_AND2</type>
<position>194.5,-74.5</position>
<input>
<ID>IN_0</ID>21 </input>
<input>
<ID>IN_1</ID>20 </input>
<output>
<ID>OUT</ID>26 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>77</ID>
<type>GA_LED</type>
<position>202.5,-74.5</position>
<input>
<ID>N_in0</ID>26 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>78</ID>
<type>AA_LABEL</type>
<position>210,-74</position>
<gparam>LABEL_TEXT BORROW(A'B)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>107,-34.5,107,-32</points>
<intersection>-34.5 1</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>107,-34.5,109.5,-34.5</points>
<connection>
<GID>55</GID>
<name>IN_0</name></connection>
<intersection>107 0</intersection>
<intersection>107.5 3</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104.5,-32,107,-32</points>
<connection>
<GID>53</GID>
<name>OUT_0</name></connection>
<intersection>107 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>107.5,-42,107.5,-34.5</points>
<intersection>-42 4</intersection>
<intersection>-34.5 1</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>107.5,-42,111,-42</points>
<connection>
<GID>57</GID>
<name>IN_0</name></connection>
<intersection>107.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106.5,-51.5,106.5,-36.5</points>
<intersection>-51.5 3</intersection>
<intersection>-39 2</intersection>
<intersection>-36.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106.5,-36.5,109.5,-36.5</points>
<connection>
<GID>55</GID>
<name>IN_1</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>104,-39,106.5,-39</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>106.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>106.5,-51.5,115,-51.5</points>
<connection>
<GID>58</GID>
<name>IN_1</name></connection>
<intersection>106.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>115.5,-35.5,117,-35.5</points>
<connection>
<GID>56</GID>
<name>N_in0</name></connection>
<connection>
<GID>55</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>111,-49.5,111,-48</points>
<connection>
<GID>57</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-49.5,115,-49.5</points>
<connection>
<GID>58</GID>
<name>IN_0</name></connection>
<intersection>111 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>121,-50.5,124.5,-50.5</points>
<connection>
<GID>59</GID>
<name>N_in0</name></connection>
<connection>
<GID>58</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>163.5,-62,163.5,-37</points>
<connection>
<GID>67</GID>
<name>OUT_0</name></connection>
<intersection>-62 3</intersection>
<intersection>-41.5 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>163.5,-62,190.5,-62</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>163.5,-41.5,170,-41.5</points>
<connection>
<GID>69</GID>
<name>IN_0</name></connection>
<intersection>163.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>20</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>175,-75.5,175,-37</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>-75.5 6</intersection>
<intersection>-55 3</intersection>
<intersection>-41 4</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>175,-55,190,-55</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>175 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>175,-41,183.5,-41</points>
<connection>
<GID>70</GID>
<name>IN_0</name></connection>
<intersection>175 0</intersection></hsegment>
<hsegment>
<ID>6</ID>
<points>175,-75.5,191.5,-75.5</points>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>175 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>170,-73.5,170,-47.5</points>
<connection>
<GID>69</GID>
<name>OUT_0</name></connection>
<intersection>-73.5 3</intersection>
<intersection>-53 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>170,-53,190,-53</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>170,-73.5,191.5,-73.5</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<intersection>170 0</intersection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>183.5,-64,183.5,-47</points>
<connection>
<GID>70</GID>
<name>OUT_0</name></connection>
<intersection>-64 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>183.5,-64,190.5,-64</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>183.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>23</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-57.5,198,-54</points>
<intersection>-57.5 2</intersection>
<intersection>-54 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196,-54,198,-54</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198,-57.5,200,-57.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>198 0</intersection></hsegment></shape></wire>
<wire>
<ID>24</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>198,-63,198,-59.5</points>
<intersection>-63 1</intersection>
<intersection>-59.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>196.5,-63,198,-63</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>198 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>198,-59.5,200,-59.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>198 0</intersection></hsegment></shape></wire>
<wire>
<ID>25</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>206,-58.5,206,-58.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<connection>
<GID>74</GID>
<name>N_in0</name></connection></vsegment></shape></wire>
<wire>
<ID>26</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>197.5,-74.5,201.5,-74.5</points>
<connection>
<GID>77</GID>
<name>N_in0</name></connection>
<connection>
<GID>76</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>44.7,-8,167.1,-68.5</PageViewport>
<gate>
<ID>1</ID>
<type>AA_LABEL</type>
<position>80.5,-17.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>2</ID>
<type>AA_LABEL</type>
<position>97,-17.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>3</ID>
<type>AA_TOGGLE</type>
<position>80.5,-21.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>97,-21.5</position>
<output>
<ID>OUT_0</ID>2 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>5</ID>
<type>BA_NAND2</type>
<position>85,-30.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>6</ID>
<type>BA_NAND2</type>
<position>102,-30</position>
<input>
<ID>IN_0</ID>2 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>7</ID>
<type>BA_NAND2</type>
<position>107.5,-45</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>5 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>BA_NAND2</type>
<position>108,-53.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>6 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>9</ID>
<type>BA_NAND2</type>
<position>117,-49</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>GA_LED</type>
<position>124,-49.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>BA_NAND2</type>
<position>108,-63</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>13</ID>
<type>BA_NAND2</type>
<position>117,-63</position>
<input>
<ID>IN_0</ID>8 </input>
<input>
<ID>IN_1</ID>8 </input>
<output>
<ID>OUT</ID>9 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>14</ID>
<type>GA_LED</type>
<position>125,-62.5</position>
<input>
<ID>N_in0</ID>9 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>AA_LABEL</type>
<position>93,-12</position>
<gparam>LABEL_TEXT NAND IMPLEMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_LABEL</type>
<position>134.5,-49</position>
<gparam>LABEL_TEXT DIFFERENCE(A'B+AB')</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0</gparam></gate>
<gate>
<ID>19</ID>
<type>AA_LABEL</type>
<position>133,-62</position>
<gparam>LABEL_TEXT BORROW(A'B)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>80.5,-27.5,86,-27.5</points>
<connection>
<GID>5</GID>
<name>IN_1</name></connection>
<connection>
<GID>5</GID>
<name>IN_0</name></connection>
<intersection>80.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>80.5,-54.5,80.5,-23.5</points>
<connection>
<GID>3</GID>
<name>OUT_0</name></connection>
<intersection>-54.5 5</intersection>
<intersection>-27.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>80.5,-54.5,105,-54.5</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>80.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>97,-27,103,-27</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<connection>
<GID>6</GID>
<name>IN_0</name></connection>
<intersection>97 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>97,-64,97,-23.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-64 9</intersection>
<intersection>-46 5</intersection>
<intersection>-27 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>97,-46,104.5,-46</points>
<connection>
<GID>7</GID>
<name>IN_1</name></connection>
<intersection>97 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>97,-64,105,-64</points>
<connection>
<GID>12</GID>
<name>IN_1</name></connection>
<intersection>97 3</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>85,-62,85,-33.5</points>
<connection>
<GID>5</GID>
<name>OUT</name></connection>
<intersection>-62 3</intersection>
<intersection>-44 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>85,-44,104.5,-44</points>
<connection>
<GID>7</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>85,-62,105,-62</points>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>85 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>102,-52.5,102,-33</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>102,-52.5,105,-52.5</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>102 0</intersection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112,-48,112,-45</points>
<intersection>-48 1</intersection>
<intersection>-45 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112,-48,114,-48</points>
<connection>
<GID>9</GID>
<name>IN_0</name></connection>
<intersection>112 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>110.5,-45,112,-45</points>
<connection>
<GID>7</GID>
<name>OUT</name></connection>
<intersection>112 0</intersection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>112.5,-53.5,112.5,-50</points>
<intersection>-53.5 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>112.5,-50,114,-50</points>
<connection>
<GID>9</GID>
<name>IN_1</name></connection>
<intersection>112.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>111,-53.5,112.5,-53.5</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>112.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>121.5,-49.5,121.5,-49</points>
<intersection>-49.5 1</intersection>
<intersection>-49 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>121.5,-49.5,123,-49.5</points>
<connection>
<GID>10</GID>
<name>N_in0</name></connection>
<intersection>121.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-49,121.5,-49</points>
<connection>
<GID>9</GID>
<name>OUT</name></connection>
<intersection>121.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>114,-64,114,-62</points>
<connection>
<GID>13</GID>
<name>IN_1</name></connection>
<connection>
<GID>13</GID>
<name>IN_0</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>111,-63,114,-63</points>
<connection>
<GID>12</GID>
<name>OUT</name></connection>
<intersection>114 0</intersection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>122,-63,122,-62.5</points>
<intersection>-63 2</intersection>
<intersection>-62.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>122,-62.5,124,-62.5</points>
<connection>
<GID>14</GID>
<name>N_in0</name></connection>
<intersection>122 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>120,-63,122,-63</points>
<connection>
<GID>13</GID>
<name>OUT</name></connection>
<intersection>122 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-17.1,7.56667,146.1,-73.1</PageViewport>
<gate>
<ID>11</ID>
<type>AA_LABEL</type>
<position>39,-2.5</position>
<gparam>LABEL_TEXT NOR IMPLEMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>15</ID>
<type>AA_LABEL</type>
<position>25,-6.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>17</ID>
<type>AA_LABEL</type>
<position>41.5,-6.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_TOGGLE</type>
<position>25,-10.5</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>41.5,-10.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>22</ID>
<type>GA_LED</type>
<position>78,-37</position>
<input>
<ID>N_in0</ID>30 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>23</ID>
<type>AA_LABEL</type>
<position>86.5,-37</position>
<gparam>LABEL_TEXT SUM[(A'B)(AB')]'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>GA_LED</type>
<position>69.5,-51.5</position>
<input>
<ID>N_in0</ID>31 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>77,-51.5</position>
<gparam>LABEL_TEXT CARRY((AB)')'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>BE_NOR2</type>
<position>31.5,-17.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>10 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>27</ID>
<type>BE_NOR2</type>
<position>47,-17</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>BE_NOR2</type>
<position>51.5,-34.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>28 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>BE_NOR2</type>
<position>52,-41</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>27 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>30</ID>
<type>BE_NOR2</type>
<position>61,-37.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>27 </input>
<output>
<ID>OUT</ID>29 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>31</ID>
<type>BE_NOR2</type>
<position>53,-51.5</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>32</ID>
<type>BE_NOR2</type>
<position>70,-37.5</position>
<input>
<ID>IN_0</ID>29 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>10</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>25,-14.5,32.5,-14.5</points>
<connection>
<GID>26</GID>
<name>IN_1</name></connection>
<connection>
<GID>26</GID>
<name>IN_0</name></connection>
<intersection>25 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>25,-50.5,25,-12.5</points>
<connection>
<GID>20</GID>
<name>OUT_0</name></connection>
<intersection>-50.5 9</intersection>
<intersection>-33.5 5</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>25,-33.5,48.5,-33.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<intersection>25 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>25,-50.5,50,-50.5</points>
<connection>
<GID>31</GID>
<name>IN_0</name></connection>
<intersection>25 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>41.5,-14,48,-14</points>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<intersection>41.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>41.5,-40,41.5,-12.5</points>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection>
<intersection>-40 5</intersection>
<intersection>-14 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>41.5,-40,49,-40</points>
<connection>
<GID>29</GID>
<name>IN_0</name></connection>
<intersection>41.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>47,-52.5,47,-20</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>-52.5 3</intersection>
<intersection>-35.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>47,-35.5,48.5,-35.5</points>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>47 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>47,-52.5,50,-52.5</points>
<connection>
<GID>31</GID>
<name>IN_1</name></connection>
<intersection>47 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>31.5,-42,31.5,-20.5</points>
<connection>
<GID>26</GID>
<name>OUT</name></connection>
<intersection>-42 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>31.5,-42,49,-42</points>
<connection>
<GID>29</GID>
<name>IN_1</name></connection>
<intersection>31.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>27</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56.5,-41,56.5,-38.5</points>
<intersection>-41 2</intersection>
<intersection>-38.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56.5,-38.5,58,-38.5</points>
<connection>
<GID>30</GID>
<name>IN_1</name></connection>
<intersection>56.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>55,-41,56.5,-41</points>
<connection>
<GID>29</GID>
<name>OUT</name></connection>
<intersection>56.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>56,-36.5,56,-34.5</points>
<intersection>-36.5 1</intersection>
<intersection>-34.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>56,-36.5,58,-36.5</points>
<connection>
<GID>30</GID>
<name>IN_0</name></connection>
<intersection>56 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>54.5,-34.5,56,-34.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>56 0</intersection></hsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67,-38.5,67,-36.5</points>
<connection>
<GID>32</GID>
<name>IN_1</name></connection>
<connection>
<GID>32</GID>
<name>IN_0</name></connection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64,-37.5,67,-37.5</points>
<connection>
<GID>30</GID>
<name>OUT</name></connection>
<intersection>67 0</intersection></hsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-37.5,75,-37</points>
<intersection>-37.5 2</intersection>
<intersection>-37 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-37,77,-37</points>
<connection>
<GID>22</GID>
<name>N_in0</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73,-37.5,75,-37.5</points>
<connection>
<GID>32</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56,-51.5,68.5,-51.5</points>
<connection>
<GID>31</GID>
<name>OUT</name></connection>
<connection>
<GID>24</GID>
<name>N_in0</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,7.5274e-007,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,7.5274e-007,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,7.5274e-007,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,7.5274e-007,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,7.5274e-007,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,7.5274e-007,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,7.5274e-007,122.4,-60.5</PageViewport></page 9></circuit>
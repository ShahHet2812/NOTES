<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>70.5078,-8.78639,233.708,-89.4534</PageViewport>
<gate>
<ID>2</ID>
<type>AA_TOGGLE</type>
<position>90.5,-35.5</position>
<output>
<ID>OUT_0</ID>4 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>104,-35.5</position>
<output>
<ID>OUT_0</ID>3 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>AA_AND2</type>
<position>118,-46.5</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>1 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>8</ID>
<type>AA_AND2</type>
<position>118,-57</position>
<input>
<ID>IN_0</ID>6 </input>
<input>
<ID>IN_1</ID>4 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>10</ID>
<type>AE_OR2</type>
<position>128.5,-51.5</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>2 </input>
<output>
<ID>OUT</ID>7 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>12</ID>
<type>AA_INVERTER</type>
<position>90.5,-42.5</position>
<input>
<ID>IN_0</ID>4 </input>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>14</ID>
<type>AA_INVERTER</type>
<position>106,-53.5</position>
<input>
<ID>IN_0</ID>3 </input>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 1</lparam></gate>
<gate>
<ID>16</ID>
<type>GA_LED</type>
<position>134.5,-51.5</position>
<input>
<ID>N_in0</ID>7 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>18</ID>
<type>AA_AND2</type>
<position>118,-70.5</position>
<input>
<ID>IN_0</ID>4 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>8 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>20</ID>
<type>GA_LED</type>
<position>126.5,-70.5</position>
<input>
<ID>N_in0</ID>8 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>124.5,-21.5</position>
<gparam>LABEL_TEXT Half Adder Circuit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_LABEL</type>
<position>139.5,-51</position>
<gparam>LABEL_TEXT A'B+AB'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>90.5,-32.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>28</ID>
<type>AA_LABEL</type>
<position>104,-32.5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>146.5,-51</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>132.5,-70.5</position>
<gparam>LABEL_TEXT CARRY(AB)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>190,-32</position>
<output>
<ID>OUT_0</ID>10 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_TOGGLE</type>
<position>190,-36</position>
<output>
<ID>OUT_0</ID>9 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>187.5,-31.5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>36</ID>
<type>AA_LABEL</type>
<position>187.5,-36</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>38</ID>
<type>AI_XOR2</type>
<position>204,-34</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>12 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>AA_AND2</type>
<position>205.5,-42</position>
<input>
<ID>IN_0</ID>10 </input>
<input>
<ID>IN_1</ID>9 </input>
<output>
<ID>OUT</ID>11 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>42</ID>
<type>GA_LED</type>
<position>210,-34</position>
<input>
<ID>N_in0</ID>12 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>GA_LED</type>
<position>211.5,-42</position>
<input>
<ID>N_in0</ID>11 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>215,-33.5</position>
<gparam>LABEL_TEXT A'B+AB'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>222,-33.5</position>
<gparam>LABEL_TEXT SUM</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>AA_LABEL</type>
<position>217.5,-42</position>
<gparam>LABEL_TEXT CARRY(AB)</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>49</ID>
<type>AA_LABEL</type>
<position>203.5,-24</position>
<gparam>LABEL_TEXT Simplyfied Circuit</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>1</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-50.5,123,-46.5</points>
<intersection>-50.5 1</intersection>
<intersection>-46.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-50.5,125.5,-50.5</points>
<connection>
<GID>10</GID>
<name>IN_0</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-46.5,123,-46.5</points>
<connection>
<GID>6</GID>
<name>OUT</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123,-57,123,-52.5</points>
<intersection>-57 2</intersection>
<intersection>-52.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123,-52.5,125.5,-52.5</points>
<connection>
<GID>10</GID>
<name>IN_1</name></connection>
<intersection>123 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>121,-57,123,-57</points>
<connection>
<GID>8</GID>
<name>OUT</name></connection>
<intersection>123 0</intersection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>104,-47.5,104,-37.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>104,-47.5,115,-47.5</points>
<connection>
<GID>6</GID>
<name>IN_1</name></connection>
<intersection>104 0</intersection>
<intersection>106 2</intersection></hsegment>
<vsegment>
<ID>2</ID>
<points>106,-71.5,106,-47.5</points>
<connection>
<GID>14</GID>
<name>IN_0</name></connection>
<intersection>-71.5 3</intersection>
<intersection>-47.5 1</intersection></vsegment>
<hsegment>
<ID>3</ID>
<points>106,-71.5,115,-71.5</points>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>106 2</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>90.5,-58,90.5,-37.5</points>
<connection>
<GID>2</GID>
<name>OUT_0</name></connection>
<connection>
<GID>12</GID>
<name>IN_0</name></connection>
<intersection>-58 2</intersection></vsegment>
<hsegment>
<ID>2</ID>
<points>90.5,-58,115,-58</points>
<connection>
<GID>8</GID>
<name>IN_1</name></connection>
<intersection>90.5 0</intersection>
<intersection>115 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>115,-69.5,115,-58</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<intersection>-58 2</intersection></vsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>90.5,-45.5,115,-45.5</points>
<connection>
<GID>12</GID>
<name>OUT_0</name></connection>
<connection>
<GID>6</GID>
<name>IN_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>106,-56.5,106,-56</points>
<connection>
<GID>14</GID>
<name>OUT_0</name></connection>
<intersection>-56 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>106,-56,115,-56</points>
<connection>
<GID>8</GID>
<name>IN_0</name></connection>
<intersection>106 0</intersection></hsegment></shape></wire>
<wire>
<ID>7</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>131.5,-51.5,133.5,-51.5</points>
<connection>
<GID>16</GID>
<name>N_in0</name></connection>
<connection>
<GID>10</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>8</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>121,-70.5,125.5,-70.5</points>
<connection>
<GID>20</GID>
<name>N_in0</name></connection>
<connection>
<GID>18</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>9</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,-43,196.5,-35</points>
<intersection>-43 4</intersection>
<intersection>-36 1</intersection>
<intersection>-35 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-36,196.5,-36</points>
<connection>
<GID>34</GID>
<name>OUT_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>196.5,-35,201,-35</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>4</ID>
<points>196.5,-43,202.5,-43</points>
<connection>
<GID>40</GID>
<name>IN_1</name></connection>
<intersection>196.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>10</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>196.5,-33,196.5,-32</points>
<intersection>-33 2</intersection>
<intersection>-32 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>192,-32,196.5,-32</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>196.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>196.5,-33,201,-33</points>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>196.5 0</intersection>
<intersection>199 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>199,-41,199,-33</points>
<intersection>-41 4</intersection>
<intersection>-33 2</intersection></vsegment>
<hsegment>
<ID>4</ID>
<points>199,-41,202.5,-41</points>
<connection>
<GID>40</GID>
<name>IN_0</name></connection>
<intersection>199 3</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>208.5,-42,210.5,-42</points>
<connection>
<GID>44</GID>
<name>N_in0</name></connection>
<connection>
<GID>40</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>207,-34,209,-34</points>
<connection>
<GID>42</GID>
<name>N_in0</name></connection>
<connection>
<GID>38</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>-20.4,10.0667,142.8,-70.6</PageViewport>
<gate>
<ID>100</ID>
<type>AA_LABEL</type>
<position>34,-5</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>101</ID>
<type>AA_LABEL</type>
<position>50.5,-5</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>102</ID>
<type>AA_TOGGLE</type>
<position>34,-9</position>
<output>
<ID>OUT_0</ID>54 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>103</ID>
<type>AA_TOGGLE</type>
<position>50.5,-9</position>
<output>
<ID>OUT_0</ID>55 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>104</ID>
<type>BA_NAND2</type>
<position>38.5,-18</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>56 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>105</ID>
<type>BA_NAND2</type>
<position>55.5,-17.5</position>
<input>
<ID>IN_0</ID>55 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>57 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>106</ID>
<type>BA_NAND2</type>
<position>61,-32.5</position>
<input>
<ID>IN_0</ID>56 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>58 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>107</ID>
<type>BA_NAND2</type>
<position>61.5,-41</position>
<input>
<ID>IN_0</ID>57 </input>
<input>
<ID>IN_1</ID>54 </input>
<output>
<ID>OUT</ID>59 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>108</ID>
<type>BA_NAND2</type>
<position>70.5,-36.5</position>
<input>
<ID>IN_0</ID>58 </input>
<input>
<ID>IN_1</ID>59 </input>
<output>
<ID>OUT</ID>60 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>109</ID>
<type>GA_LED</type>
<position>77.5,-37</position>
<input>
<ID>N_in0</ID>60 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>110</ID>
<type>AA_LABEL</type>
<position>86,-37</position>
<gparam>LABEL_TEXT SUM[(A'B)(AB')]'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>111</ID>
<type>BA_NAND2</type>
<position>61.5,-50.5</position>
<input>
<ID>IN_0</ID>54 </input>
<input>
<ID>IN_1</ID>55 </input>
<output>
<ID>OUT</ID>61 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>113</ID>
<type>BA_NAND2</type>
<position>70.5,-50.5</position>
<input>
<ID>IN_0</ID>61 </input>
<input>
<ID>IN_1</ID>61 </input>
<output>
<ID>OUT</ID>62 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>115</ID>
<type>GA_LED</type>
<position>78.5,-50</position>
<input>
<ID>N_in0</ID>62 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>117</ID>
<type>AA_LABEL</type>
<position>86,-50</position>
<gparam>LABEL_TEXT CARRY((AB)')'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>119</ID>
<type>AA_LABEL</type>
<position>46.5,0.5</position>
<gparam>LABEL_TEXT NAND IMPLEMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<wire>
<ID>54</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>34,-15,39.5,-15</points>
<connection>
<GID>104</GID>
<name>IN_1</name></connection>
<connection>
<GID>104</GID>
<name>IN_0</name></connection>
<intersection>34 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>34,-49.5,34,-11</points>
<connection>
<GID>102</GID>
<name>OUT_0</name></connection>
<intersection>-49.5 9</intersection>
<intersection>-42 5</intersection>
<intersection>-15 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>34,-42,58.5,-42</points>
<connection>
<GID>107</GID>
<name>IN_1</name></connection>
<intersection>34 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>34,-49.5,58.5,-49.5</points>
<connection>
<GID>111</GID>
<name>IN_0</name></connection>
<intersection>34 3</intersection></hsegment></shape></wire>
<wire>
<ID>55</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>50.5,-14.5,56.5,-14.5</points>
<connection>
<GID>105</GID>
<name>IN_1</name></connection>
<connection>
<GID>105</GID>
<name>IN_0</name></connection>
<intersection>50.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>50.5,-51.5,50.5,-11</points>
<connection>
<GID>103</GID>
<name>OUT_0</name></connection>
<intersection>-51.5 9</intersection>
<intersection>-33.5 5</intersection>
<intersection>-14.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>50.5,-33.5,58,-33.5</points>
<connection>
<GID>106</GID>
<name>IN_1</name></connection>
<intersection>50.5 3</intersection></hsegment>
<hsegment>
<ID>9</ID>
<points>50.5,-51.5,58.5,-51.5</points>
<connection>
<GID>111</GID>
<name>IN_1</name></connection>
<intersection>50.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>56</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>38.5,-31.5,38.5,-21</points>
<connection>
<GID>104</GID>
<name>OUT</name></connection>
<intersection>-31.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>38.5,-31.5,58,-31.5</points>
<connection>
<GID>106</GID>
<name>IN_0</name></connection>
<intersection>38.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>57</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55.5,-40,55.5,-20.5</points>
<connection>
<GID>105</GID>
<name>OUT</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55.5,-40,58.5,-40</points>
<connection>
<GID>107</GID>
<name>IN_0</name></connection>
<intersection>55.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>58</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>65.5,-35.5,65.5,-32.5</points>
<intersection>-35.5 1</intersection>
<intersection>-32.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>65.5,-35.5,67.5,-35.5</points>
<connection>
<GID>108</GID>
<name>IN_0</name></connection>
<intersection>65.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64,-32.5,65.5,-32.5</points>
<connection>
<GID>106</GID>
<name>OUT</name></connection>
<intersection>65.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>59</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>66,-41,66,-37.5</points>
<intersection>-41 2</intersection>
<intersection>-37.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>66,-37.5,67.5,-37.5</points>
<connection>
<GID>108</GID>
<name>IN_1</name></connection>
<intersection>66 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>64.5,-41,66,-41</points>
<connection>
<GID>107</GID>
<name>OUT</name></connection>
<intersection>66 0</intersection></hsegment></shape></wire>
<wire>
<ID>60</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75,-37,75,-36.5</points>
<intersection>-37 1</intersection>
<intersection>-36.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75,-37,76.5,-37</points>
<connection>
<GID>109</GID>
<name>N_in0</name></connection>
<intersection>75 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-36.5,75,-36.5</points>
<connection>
<GID>108</GID>
<name>OUT</name></connection>
<intersection>75 0</intersection></hsegment></shape></wire>
<wire>
<ID>61</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>67.5,-51.5,67.5,-49.5</points>
<connection>
<GID>113</GID>
<name>IN_0</name></connection>
<connection>
<GID>113</GID>
<name>IN_1</name></connection>
<intersection>-50.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>64.5,-50.5,67.5,-50.5</points>
<connection>
<GID>111</GID>
<name>OUT</name></connection>
<intersection>67.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>62</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>75.5,-50.5,75.5,-50</points>
<intersection>-50.5 2</intersection>
<intersection>-50 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>75.5,-50,77.5,-50</points>
<connection>
<GID>115</GID>
<name>N_in0</name></connection>
<intersection>75.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>73.5,-50.5,75.5,-50.5</points>
<connection>
<GID>113</GID>
<name>OUT</name></connection>
<intersection>75.5 0</intersection></hsegment></shape></wire></page 1>
<page 2>
<PageViewport>-17.1,7.56667,146.1,-73.1</PageViewport>
<gate>
<ID>121</ID>
<type>AA_LABEL</type>
<position>52,-5</position>
<gparam>LABEL_TEXT NOR IMPLEMENTATION</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>122</ID>
<type>AA_LABEL</type>
<position>38,-9</position>
<gparam>LABEL_TEXT A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>123</ID>
<type>AA_LABEL</type>
<position>54.5,-9</position>
<gparam>LABEL_TEXT B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>124</ID>
<type>AA_TOGGLE</type>
<position>38,-13</position>
<output>
<ID>OUT_0</ID>72 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>125</ID>
<type>AA_TOGGLE</type>
<position>54.5,-13</position>
<output>
<ID>OUT_0</ID>73 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 270</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>131</ID>
<type>GA_LED</type>
<position>91,-39.5</position>
<input>
<ID>N_in0</ID>80 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>132</ID>
<type>AA_LABEL</type>
<position>99.5,-39.5</position>
<gparam>LABEL_TEXT SUM[(A'B)(AB')]'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>135</ID>
<type>GA_LED</type>
<position>82.5,-54</position>
<input>
<ID>N_in0</ID>81 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>136</ID>
<type>AA_LABEL</type>
<position>90,-54</position>
<gparam>LABEL_TEXT CARRY((AB)')'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>138</ID>
<type>BE_NOR2</type>
<position>44.5,-20</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>72 </input>
<output>
<ID>OUT</ID>75 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>140</ID>
<type>BE_NOR2</type>
<position>60,-19.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>73 </input>
<output>
<ID>OUT</ID>74 </output>
<gparam>angle 270</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>142</ID>
<type>BE_NOR2</type>
<position>64.5,-37</position>
<input>
<ID>IN_0</ID>72 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>77 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>144</ID>
<type>BE_NOR2</type>
<position>65,-43.5</position>
<input>
<ID>IN_0</ID>73 </input>
<input>
<ID>IN_1</ID>75 </input>
<output>
<ID>OUT</ID>76 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>148</ID>
<type>BE_NOR2</type>
<position>74,-40</position>
<input>
<ID>IN_0</ID>77 </input>
<input>
<ID>IN_1</ID>76 </input>
<output>
<ID>OUT</ID>79 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>152</ID>
<type>BE_NOR2</type>
<position>66,-54</position>
<input>
<ID>IN_0</ID>75 </input>
<input>
<ID>IN_1</ID>74 </input>
<output>
<ID>OUT</ID>81 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>156</ID>
<type>BE_NOR2</type>
<position>83,-40</position>
<input>
<ID>IN_0</ID>79 </input>
<input>
<ID>IN_1</ID>79 </input>
<output>
<ID>OUT</ID>80 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>72</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>38,-17,45.5,-17</points>
<connection>
<GID>138</GID>
<name>IN_0</name></connection>
<connection>
<GID>138</GID>
<name>IN_1</name></connection>
<intersection>38 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>38,-36,38,-15</points>
<connection>
<GID>124</GID>
<name>OUT_0</name></connection>
<intersection>-36 5</intersection>
<intersection>-17 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>38,-36,61.5,-36</points>
<connection>
<GID>142</GID>
<name>IN_0</name></connection>
<intersection>38 3</intersection></hsegment></shape></wire>
<wire>
<ID>73</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>54.5,-16.5,61,-16.5</points>
<connection>
<GID>140</GID>
<name>IN_0</name></connection>
<connection>
<GID>140</GID>
<name>IN_1</name></connection>
<intersection>54.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>54.5,-42.5,54.5,-15</points>
<connection>
<GID>125</GID>
<name>OUT_0</name></connection>
<intersection>-42.5 5</intersection>
<intersection>-16.5 1</intersection></vsegment>
<hsegment>
<ID>5</ID>
<points>54.5,-42.5,62,-42.5</points>
<connection>
<GID>144</GID>
<name>IN_0</name></connection>
<intersection>54.5 3</intersection></hsegment></shape></wire>
<wire>
<ID>74</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>60,-55,60,-22.5</points>
<connection>
<GID>140</GID>
<name>OUT</name></connection>
<intersection>-55 3</intersection>
<intersection>-38 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>60,-38,61.5,-38</points>
<connection>
<GID>142</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>60,-55,63,-55</points>
<connection>
<GID>152</GID>
<name>IN_1</name></connection>
<intersection>60 0</intersection></hsegment></shape></wire>
<wire>
<ID>75</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>44.5,-53,44.5,-23</points>
<connection>
<GID>138</GID>
<name>OUT</name></connection>
<intersection>-53 3</intersection>
<intersection>-44.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>44.5,-44.5,62,-44.5</points>
<connection>
<GID>144</GID>
<name>IN_1</name></connection>
<intersection>44.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>44.5,-53,63,-53</points>
<connection>
<GID>152</GID>
<name>IN_0</name></connection>
<intersection>44.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>76</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69.5,-43.5,69.5,-41</points>
<intersection>-43.5 2</intersection>
<intersection>-41 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69.5,-41,71,-41</points>
<connection>
<GID>148</GID>
<name>IN_1</name></connection>
<intersection>69.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>68,-43.5,69.5,-43.5</points>
<connection>
<GID>144</GID>
<name>OUT</name></connection>
<intersection>69.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>77</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>69,-39,69,-37</points>
<intersection>-39 1</intersection>
<intersection>-37 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>69,-39,71,-39</points>
<connection>
<GID>148</GID>
<name>IN_0</name></connection>
<intersection>69 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>67.5,-37,69,-37</points>
<connection>
<GID>142</GID>
<name>OUT</name></connection>
<intersection>69 0</intersection></hsegment></shape></wire>
<wire>
<ID>79</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>80,-41,80,-39</points>
<connection>
<GID>156</GID>
<name>IN_0</name></connection>
<connection>
<GID>156</GID>
<name>IN_1</name></connection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>77,-40,80,-40</points>
<connection>
<GID>148</GID>
<name>OUT</name></connection>
<intersection>80 0</intersection></hsegment></shape></wire>
<wire>
<ID>80</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>88,-40,88,-39.5</points>
<intersection>-40 2</intersection>
<intersection>-39.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>88,-39.5,90,-39.5</points>
<connection>
<GID>131</GID>
<name>N_in0</name></connection>
<intersection>88 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>86,-40,88,-40</points>
<connection>
<GID>156</GID>
<name>OUT</name></connection>
<intersection>88 0</intersection></hsegment></shape></wire>
<wire>
<ID>81</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>69,-54,81.5,-54</points>
<connection>
<GID>135</GID>
<name>N_in0</name></connection>
<connection>
<GID>152</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 2>
<page 3>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,7.42428e-007,122.4,-60.5</PageViewport></page 9></circuit>
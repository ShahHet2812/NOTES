<circuit>
<CurrentPage>0</CurrentPage>
<page 0>
<PageViewport>-12.2918,0.369435,205.308,-107.186</PageViewport>
<gate>
<ID>2</ID>
<type>BA_NAND2</type>
<position>45,-25</position>
<input>
<ID>IN_0</ID>1 </input>
<input>
<ID>IN_1</ID>1 </input>
<output>
<ID>OUT</ID>2 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>4</ID>
<type>AA_TOGGLE</type>
<position>30.5,-25.5</position>
<output>
<ID>OUT_0</ID>1 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>6</ID>
<type>GA_LED</type>
<position>53,-25</position>
<input>
<ID>N_in0</ID>2 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>8</ID>
<type>AA_LABEL</type>
<position>24,-25</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>10</ID>
<type>AA_LABEL</type>
<position>60,-24.5</position>
<gparam>LABEL_TEXT Output Y=A'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>12</ID>
<type>AA_LABEL</type>
<position>44.5,-18</position>
<gparam>LABEL_TEXT NAND as NOT Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>14</ID>
<type>AA_LABEL</type>
<position>93.5,-7.5</position>
<gparam>LABEL_TEXT NAND Gate as UNIVERSAL GATE</gparam>
<gparam>TEXT_HEIGHT 3</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>16</ID>
<type>BA_NAND2</type>
<position>39,-39</position>
<input>
<ID>IN_0</ID>5 </input>
<input>
<ID>IN_1</ID>6 </input>
<output>
<ID>OUT</ID>3 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>18</ID>
<type>BA_NAND2</type>
<position>53.5,-39</position>
<input>
<ID>IN_0</ID>3 </input>
<input>
<ID>IN_1</ID>3 </input>
<output>
<ID>OUT</ID>4 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>19</ID>
<type>GA_LED</type>
<position>60.5,-39</position>
<input>
<ID>N_in0</ID>4 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>20</ID>
<type>AA_LABEL</type>
<position>67.5,-38.5</position>
<gparam>LABEL_TEXT Output Y=A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>21</ID>
<type>AA_TOGGLE</type>
<position>29,-38</position>
<output>
<ID>OUT_0</ID>5 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 1</lparam></gate>
<gate>
<ID>22</ID>
<type>AA_LABEL</type>
<position>22.5,-37.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>24</ID>
<type>AA_TOGGLE</type>
<position>29,-41</position>
<output>
<ID>OUT_0</ID>6 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>25</ID>
<type>AA_LABEL</type>
<position>23,-41</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>26</ID>
<type>AA_LABEL</type>
<position>45,-32.5</position>
<gparam>LABEL_TEXT NAND as AND Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>27</ID>
<type>BA_NAND2</type>
<position>38,-58.5</position>
<input>
<ID>IN_0</ID>11 </input>
<input>
<ID>IN_1</ID>11 </input>
<output>
<ID>OUT</ID>14 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>28</ID>
<type>BA_NAND2</type>
<position>38,-65.5</position>
<input>
<ID>IN_0</ID>12 </input>
<input>
<ID>IN_1</ID>12 </input>
<output>
<ID>OUT</ID>13 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>29</ID>
<type>GA_LED</type>
<position>59.5,-58.5</position>
<input>
<ID>N_in0</ID>15 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>30</ID>
<type>AA_LABEL</type>
<position>66.5,-58</position>
<gparam>LABEL_TEXT Output Y=A.B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>31</ID>
<type>AA_TOGGLE</type>
<position>28,-57.5</position>
<output>
<ID>OUT_0</ID>11 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>32</ID>
<type>AA_LABEL</type>
<position>21.5,-57</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>33</ID>
<type>AA_TOGGLE</type>
<position>28,-66</position>
<output>
<ID>OUT_0</ID>12 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>34</ID>
<type>AA_LABEL</type>
<position>22.5,-66</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>35</ID>
<type>AA_LABEL</type>
<position>45,-50.5</position>
<gparam>LABEL_TEXT NAND as OR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>37</ID>
<type>BA_NAND2</type>
<position>49,-61</position>
<input>
<ID>IN_0</ID>14 </input>
<input>
<ID>IN_1</ID>13 </input>
<output>
<ID>OUT</ID>15 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>38</ID>
<type>BA_NAND2</type>
<position>36,-83</position>
<input>
<ID>IN_0</ID>16 </input>
<input>
<ID>IN_1</ID>16 </input>
<output>
<ID>OUT</ID>19 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>39</ID>
<type>BA_NAND2</type>
<position>36,-90</position>
<input>
<ID>IN_0</ID>17 </input>
<input>
<ID>IN_1</ID>17 </input>
<output>
<ID>OUT</ID>18 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>40</ID>
<type>GA_LED</type>
<position>59,-85.5</position>
<input>
<ID>N_in0</ID>21 </input>
<input>
<ID>N_in1</ID>21 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>41</ID>
<type>AA_LABEL</type>
<position>72.5,-85</position>
<gparam>LABEL_TEXT Output Y=(A+B)'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>42</ID>
<type>AA_TOGGLE</type>
<position>26,-82</position>
<output>
<ID>OUT_0</ID>16 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>43</ID>
<type>AA_LABEL</type>
<position>19.5,-81.5</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>44</ID>
<type>AA_TOGGLE</type>
<position>26,-90.5</position>
<output>
<ID>OUT_0</ID>17 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>45</ID>
<type>AA_LABEL</type>
<position>20.5,-90.5</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>46</ID>
<type>AA_LABEL</type>
<position>43,-75</position>
<gparam>LABEL_TEXT NAND as NOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>47</ID>
<type>BA_NAND2</type>
<position>47,-85.5</position>
<input>
<ID>IN_0</ID>19 </input>
<input>
<ID>IN_1</ID>18 </input>
<output>
<ID>OUT</ID>22 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>49</ID>
<type>BA_NAND2</type>
<position>54,-85.5</position>
<input>
<ID>IN_0</ID>22 </input>
<input>
<ID>IN_1</ID>22 </input>
<output>
<ID>OUT</ID>21 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>52</ID>
<type>GA_LED</type>
<position>146,-24.5</position>
<input>
<ID>N_in0</ID>33 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>53</ID>
<type>AA_LABEL</type>
<position>155,-24</position>
<gparam>LABEL_TEXT Output Y=A'B+AB'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>54</ID>
<type>AA_TOGGLE</type>
<position>114.5,-23.5</position>
<output>
<ID>OUT_0</ID>28 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>55</ID>
<type>AA_LABEL</type>
<position>108,-23</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>56</ID>
<type>AA_TOGGLE</type>
<position>114.5,-32</position>
<output>
<ID>OUT_0</ID>29 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>57</ID>
<type>AA_LABEL</type>
<position>109,-32</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>58</ID>
<type>AA_LABEL</type>
<position>131.5,-16.5</position>
<gparam>LABEL_TEXT NAND as XOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>59</ID>
<type>BA_NAND2</type>
<position>124.5,-27.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>30 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>60</ID>
<type>BA_NAND2</type>
<position>134.5,-23.5</position>
<input>
<ID>IN_0</ID>28 </input>
<input>
<ID>IN_1</ID>30 </input>
<output>
<ID>OUT</ID>31 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>61</ID>
<type>BA_NAND2</type>
<position>134,-31.5</position>
<input>
<ID>IN_0</ID>30 </input>
<input>
<ID>IN_1</ID>29 </input>
<output>
<ID>OUT</ID>32 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>63</ID>
<type>BA_NAND2</type>
<position>141,-27</position>
<input>
<ID>IN_0</ID>31 </input>
<input>
<ID>IN_1</ID>32 </input>
<output>
<ID>OUT</ID>33 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>64</ID>
<type>GA_LED</type>
<position>157.5,-64</position>
<input>
<ID>N_in0</ID>41 </input>
<gparam>LED_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>65</ID>
<type>AA_LABEL</type>
<position>166.5,-63.5</position>
<gparam>LABEL_TEXT Output Y=A'B+AB'</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>66</ID>
<type>AA_TOGGLE</type>
<position>115,-60.5</position>
<output>
<ID>OUT_0</ID>34 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>67</ID>
<type>AA_LABEL</type>
<position>108.5,-60</position>
<gparam>LABEL_TEXT Input A</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>68</ID>
<type>AA_TOGGLE</type>
<position>115,-69</position>
<output>
<ID>OUT_0</ID>35 </output>
<gparam>CLICK_BOX -0.76,-0.76,0.76,0.76</gparam>
<gparam>angle 0.0</gparam>
<lparam>OUTPUT_BITS 1</lparam>
<lparam>OUTPUT_NUM 0</lparam></gate>
<gate>
<ID>69</ID>
<type>AA_LABEL</type>
<position>109.5,-69</position>
<gparam>LABEL_TEXT Input B</gparam>
<gparam>TEXT_HEIGHT 1</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>70</ID>
<type>AA_LABEL</type>
<position>132,-53.5</position>
<gparam>LABEL_TEXT NAND as XNOR Gate</gparam>
<gparam>TEXT_HEIGHT 2</gparam>
<gparam>angle 0.0</gparam></gate>
<gate>
<ID>71</ID>
<type>BA_NAND2</type>
<position>125,-64.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>36 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>72</ID>
<type>BA_NAND2</type>
<position>135,-60.5</position>
<input>
<ID>IN_0</ID>34 </input>
<input>
<ID>IN_1</ID>36 </input>
<output>
<ID>OUT</ID>37 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>73</ID>
<type>BA_NAND2</type>
<position>134.5,-68.5</position>
<input>
<ID>IN_0</ID>36 </input>
<input>
<ID>IN_1</ID>35 </input>
<output>
<ID>OUT</ID>38 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>74</ID>
<type>BA_NAND2</type>
<position>141.5,-64</position>
<input>
<ID>IN_0</ID>37 </input>
<input>
<ID>IN_1</ID>38 </input>
<output>
<ID>OUT</ID>40 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<gate>
<ID>76</ID>
<type>BA_NAND2</type>
<position>149.5,-64</position>
<input>
<ID>IN_0</ID>40 </input>
<input>
<ID>IN_1</ID>40 </input>
<output>
<ID>OUT</ID>41 </output>
<gparam>angle 0.0</gparam>
<lparam>INPUT_BITS 2</lparam></gate>
<wire>
<ID>1</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>32.5,-25.5,42,-25.5</points>
<connection>
<GID>4</GID>
<name>OUT_0</name></connection>
<intersection>42 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>42,-26,42,-24</points>
<connection>
<GID>2</GID>
<name>IN_1</name></connection>
<connection>
<GID>2</GID>
<name>IN_0</name></connection>
<intersection>-25.5 1</intersection></vsegment></shape></wire>
<wire>
<ID>2</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>48,-25,52,-25</points>
<connection>
<GID>2</GID>
<name>OUT</name></connection>
<connection>
<GID>6</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>3</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>50.5,-40,50.5,-38</points>
<connection>
<GID>18</GID>
<name>IN_0</name></connection>
<connection>
<GID>18</GID>
<name>IN_1</name></connection>
<intersection>-39 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>42,-39,50.5,-39</points>
<connection>
<GID>16</GID>
<name>OUT</name></connection>
<intersection>50.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>4</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>56.5,-39,59.5,-39</points>
<connection>
<GID>19</GID>
<name>N_in0</name></connection>
<connection>
<GID>18</GID>
<name>OUT</name></connection></hsegment></shape></wire>
<wire>
<ID>5</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>31,-38,36,-38</points>
<connection>
<GID>16</GID>
<name>IN_0</name></connection>
<connection>
<GID>21</GID>
<name>OUT_0</name></connection></hsegment></shape></wire>
<wire>
<ID>6</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33.5,-41,33.5,-40</points>
<intersection>-41 2</intersection>
<intersection>-40 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>33.5,-40,36,-40</points>
<connection>
<GID>16</GID>
<name>IN_1</name></connection>
<intersection>33.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>31,-41,33.5,-41</points>
<connection>
<GID>24</GID>
<name>OUT_0</name></connection>
<intersection>33.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>11</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-59.5,35,-57.5</points>
<connection>
<GID>27</GID>
<name>IN_0</name></connection>
<connection>
<GID>27</GID>
<name>IN_1</name></connection>
<intersection>-57.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-57.5,35,-57.5</points>
<connection>
<GID>31</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>12</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>35,-66.5,35,-64.5</points>
<connection>
<GID>28</GID>
<name>IN_0</name></connection>
<connection>
<GID>28</GID>
<name>IN_1</name></connection>
<intersection>-66 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>30,-66,35,-66</points>
<connection>
<GID>33</GID>
<name>OUT_0</name></connection>
<intersection>35 0</intersection></hsegment></shape></wire>
<wire>
<ID>13</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-65.5,43.5,-62</points>
<intersection>-65.5 2</intersection>
<intersection>-62 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-62,46,-62</points>
<connection>
<GID>37</GID>
<name>IN_1</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-65.5,43.5,-65.5</points>
<connection>
<GID>28</GID>
<name>OUT</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>14</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>43.5,-60,43.5,-58.5</points>
<intersection>-60 1</intersection>
<intersection>-58.5 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>43.5,-60,46,-60</points>
<connection>
<GID>37</GID>
<name>IN_0</name></connection>
<intersection>43.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>41,-58.5,43.5,-58.5</points>
<connection>
<GID>27</GID>
<name>OUT</name></connection>
<intersection>43.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>15</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>55,-61,55,-58.5</points>
<intersection>-61 2</intersection>
<intersection>-58.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>55,-58.5,58.5,-58.5</points>
<connection>
<GID>29</GID>
<name>N_in0</name></connection>
<intersection>55 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>52,-61,55,-61</points>
<connection>
<GID>37</GID>
<name>OUT</name></connection>
<intersection>55 0</intersection></hsegment></shape></wire>
<wire>
<ID>16</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-84,33,-82</points>
<connection>
<GID>38</GID>
<name>IN_1</name></connection>
<connection>
<GID>38</GID>
<name>IN_0</name></connection>
<intersection>-82 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-82,33,-82</points>
<connection>
<GID>42</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>17</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>33,-91,33,-89</points>
<connection>
<GID>39</GID>
<name>IN_1</name></connection>
<connection>
<GID>39</GID>
<name>IN_0</name></connection>
<intersection>-90.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>28,-90.5,33,-90.5</points>
<connection>
<GID>44</GID>
<name>OUT_0</name></connection>
<intersection>33 0</intersection></hsegment></shape></wire>
<wire>
<ID>18</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-90,41.5,-86.5</points>
<intersection>-90 2</intersection>
<intersection>-86.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-86.5,44,-86.5</points>
<connection>
<GID>47</GID>
<name>IN_1</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-90,41.5,-90</points>
<connection>
<GID>39</GID>
<name>OUT</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>19</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>41.5,-84.5,41.5,-83</points>
<intersection>-84.5 1</intersection>
<intersection>-83 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>41.5,-84.5,44,-84.5</points>
<connection>
<GID>47</GID>
<name>IN_0</name></connection>
<intersection>41.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>39,-83,41.5,-83</points>
<connection>
<GID>38</GID>
<name>OUT</name></connection>
<intersection>41.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>21</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>57,-85.5,60,-85.5</points>
<connection>
<GID>49</GID>
<name>OUT</name></connection>
<connection>
<GID>40</GID>
<name>N_in1</name></connection>
<connection>
<GID>40</GID>
<name>N_in0</name></connection></hsegment></shape></wire>
<wire>
<ID>22</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>51,-86.5,51,-84.5</points>
<connection>
<GID>49</GID>
<name>IN_0</name></connection>
<connection>
<GID>49</GID>
<name>IN_1</name></connection>
<intersection>-85.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>50,-85.5,51,-85.5</points>
<connection>
<GID>47</GID>
<name>OUT</name></connection>
<intersection>51 0</intersection></hsegment></shape></wire>
<wire>
<ID>28</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-23.5,124,-22.5</points>
<intersection>-23.5 2</intersection>
<intersection>-22.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,-22.5,131.5,-22.5</points>
<connection>
<GID>60</GID>
<name>IN_0</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-23.5,124,-23.5</points>
<connection>
<GID>54</GID>
<name>OUT_0</name></connection>
<intersection>121.5 3</intersection>
<intersection>124 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>121.5,-26.5,121.5,-23.5</points>
<connection>
<GID>59</GID>
<name>IN_0</name></connection>
<intersection>-23.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>29</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>123.5,-32.5,123.5,-32</points>
<intersection>-32.5 1</intersection>
<intersection>-32 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>123.5,-32.5,131,-32.5</points>
<connection>
<GID>61</GID>
<name>IN_1</name></connection>
<intersection>123.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>116.5,-32,123.5,-32</points>
<connection>
<GID>56</GID>
<name>OUT_0</name></connection>
<intersection>121.5 3</intersection>
<intersection>123.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>121.5,-32,121.5,-28.5</points>
<connection>
<GID>59</GID>
<name>IN_1</name></connection>
<intersection>-32 2</intersection></vsegment></shape></wire>
<wire>
<ID>30</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129,-30.5,129,-24.5</points>
<intersection>-30.5 1</intersection>
<intersection>-27.5 2</intersection>
<intersection>-24.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129,-30.5,131,-30.5</points>
<connection>
<GID>61</GID>
<name>IN_0</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>127.5,-27.5,129,-27.5</points>
<connection>
<GID>59</GID>
<name>OUT</name></connection>
<intersection>129 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>129,-24.5,131.5,-24.5</points>
<connection>
<GID>60</GID>
<name>IN_1</name></connection>
<intersection>129 0</intersection></hsegment></shape></wire>
<wire>
<ID>31</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-26,137.5,-23.5</points>
<connection>
<GID>60</GID>
<name>OUT</name></connection>
<intersection>-26 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,-26,138,-26</points>
<connection>
<GID>63</GID>
<name>IN_0</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>32</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>137.5,-31.5,137.5,-28</points>
<intersection>-31.5 2</intersection>
<intersection>-28 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>137.5,-28,138,-28</points>
<connection>
<GID>63</GID>
<name>IN_1</name></connection>
<intersection>137.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137,-31.5,137.5,-31.5</points>
<connection>
<GID>61</GID>
<name>OUT</name></connection>
<intersection>137.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>33</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>144.5,-27,144.5,-24.5</points>
<intersection>-27 2</intersection>
<intersection>-24.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>144.5,-24.5,145,-24.5</points>
<connection>
<GID>52</GID>
<name>N_in0</name></connection>
<intersection>144.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>144,-27,144.5,-27</points>
<connection>
<GID>63</GID>
<name>OUT</name></connection>
<intersection>144.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>34</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124.5,-60.5,124.5,-59.5</points>
<intersection>-60.5 2</intersection>
<intersection>-59.5 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124.5,-59.5,132,-59.5</points>
<connection>
<GID>72</GID>
<name>IN_0</name></connection>
<intersection>124.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117,-60.5,124.5,-60.5</points>
<connection>
<GID>66</GID>
<name>OUT_0</name></connection>
<intersection>122 3</intersection>
<intersection>124.5 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>122,-63.5,122,-60.5</points>
<connection>
<GID>71</GID>
<name>IN_0</name></connection>
<intersection>-60.5 2</intersection></vsegment></shape></wire>
<wire>
<ID>35</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>124,-69.5,124,-69</points>
<intersection>-69.5 1</intersection>
<intersection>-69 2</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>124,-69.5,131.5,-69.5</points>
<connection>
<GID>73</GID>
<name>IN_1</name></connection>
<intersection>124 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>117,-69,124,-69</points>
<connection>
<GID>68</GID>
<name>OUT_0</name></connection>
<intersection>122 3</intersection>
<intersection>124 0</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>122,-69,122,-65.5</points>
<connection>
<GID>71</GID>
<name>IN_1</name></connection>
<intersection>-69 2</intersection></vsegment></shape></wire>
<wire>
<ID>36</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>129.5,-67.5,129.5,-61.5</points>
<intersection>-67.5 1</intersection>
<intersection>-64.5 2</intersection>
<intersection>-61.5 3</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>129.5,-67.5,131.5,-67.5</points>
<connection>
<GID>73</GID>
<name>IN_0</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>128,-64.5,129.5,-64.5</points>
<connection>
<GID>71</GID>
<name>OUT</name></connection>
<intersection>129.5 0</intersection></hsegment>
<hsegment>
<ID>3</ID>
<points>129.5,-61.5,132,-61.5</points>
<connection>
<GID>72</GID>
<name>IN_1</name></connection>
<intersection>129.5 0</intersection></hsegment></shape></wire>
<wire>
<ID>37</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-63,138,-60.5</points>
<connection>
<GID>72</GID>
<name>OUT</name></connection>
<intersection>-63 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-63,138.5,-63</points>
<connection>
<GID>74</GID>
<name>IN_0</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>38</ID>
<shape>
<vsegment>
<ID>0</ID>
<points>138,-68.5,138,-65</points>
<intersection>-68.5 2</intersection>
<intersection>-65 1</intersection></vsegment>
<hsegment>
<ID>1</ID>
<points>138,-65,138.5,-65</points>
<connection>
<GID>74</GID>
<name>IN_1</name></connection>
<intersection>138 0</intersection></hsegment>
<hsegment>
<ID>2</ID>
<points>137.5,-68.5,138,-68.5</points>
<connection>
<GID>73</GID>
<name>OUT</name></connection>
<intersection>138 0</intersection></hsegment></shape></wire>
<wire>
<ID>40</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>144.5,-64,146.5,-64</points>
<connection>
<GID>74</GID>
<name>OUT</name></connection>
<intersection>146.5 3</intersection>
<intersection>146.5 3</intersection></hsegment>
<vsegment>
<ID>3</ID>
<points>146.5,-65,146.5,-63</points>
<connection>
<GID>76</GID>
<name>IN_0</name></connection>
<connection>
<GID>76</GID>
<name>IN_1</name></connection>
<intersection>-64 1</intersection></vsegment></shape></wire>
<wire>
<ID>41</ID>
<shape>
<hsegment>
<ID>1</ID>
<points>152.5,-64,156.5,-64</points>
<connection>
<GID>64</GID>
<name>N_in0</name></connection>
<connection>
<GID>76</GID>
<name>OUT</name></connection></hsegment></shape></wire></page 0>
<page 1>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 1>
<page 2>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 2>
<page 3>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 3>
<page 4>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 4>
<page 5>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 5>
<page 6>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 6>
<page 7>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 7>
<page 8>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 8>
<page 9>
<PageViewport>0,3.77107e-007,122.4,-60.5</PageViewport></page 9></circuit>